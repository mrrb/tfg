/*
 * Header file for the FIFO_REG module.
 */

`ifndef _FIFO_REG_H_
`define _FIFO_REG_H_ 1

`include "FIFO_REG/rtl/FIFO_REG.v" // Main module include 

`endif