/*
 * Header file for the ULPI_REG_WRITE module.
 */

`ifndef _ULPI_REG_WRITE_H_
`define _ULPI_REG_WRITE_H_ 1

`include "ULPI/rtl/ULPI_REG_WRITE.v" // Main module include 

`endif