/*
 * Header file for the UART_Tx module.
 */

`ifndef _UART_TX_H_
`define _UART_TX_H_ 1

`include "UART/rtl/UART_Tx.v" // Main module include 

`endif