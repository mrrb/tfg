/*
 * Header file for the FIFO_BRAM_SYNC_CUSTOM module.
 */

`ifndef _FIFO_BRAM_SYNC_CUSTOM_H_
`define _FIFO_BRAM_SYNC_CUSTOM_H_ 1

`include "FIFO_BRAM_SYNC_CUSTOM/rtl/FIFO_BRAM_SYNC_CUSTOM.v" // Main module include 

`endif