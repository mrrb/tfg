/*
 * Header file for the mux module.
 */

`ifndef _MUX_H_
`define _MUX_H_ 1

`include "mux/rtl/mux.v" // Main module include 

`endif