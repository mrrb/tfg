/*
 * Header file for the ULPI_RECV module.
 */

`ifndef _ULPI_RECV_H_
`define _ULPI_RECV_H_ 1

`include "ULPI/rtl/ULPI_RECV.v" // Main module include 

`endif