/*
 * Header file for the SPI_COMM module.
 */

`ifndef _SPI_COMM_old_H_
`define _SPI_COMM_old_H_ 1

`include "SPI_COMM_old/rtl/SPI_COMM.v" // Main module include 

`endif