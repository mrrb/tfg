/*
 * Header file for the ULPI_WRAPPER module.
 */

`ifndef _ULPI_WRAPPER_H_
`define _ULPI_WRAPPER_H_ 1

`include "ULPI_WRAPPER/rtl/ULPI_WRAPPER.v" // Main module include 

`endif