/*
 * Header file for the ULPI_op_stack module.
 */

`ifndef _ULPI_OP_STACK_H_
`define _ULPI_OP_STACK_H_ 1

`include "ULPI_op_stack/rtl/ULPI_op_stack.v" // Main module include 

`endif