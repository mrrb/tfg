//! BROKEN MODULE, NOT USE!

/*
 * Header file for the FIFO_MERGE module.
 */

`ifndef _FIFO_MERGE_H_
`define _FIFO_MERGE_H_ 1

`include "FIFO_MERGE/rtl/FIFO_MERGE.v" // Main module include 

`endif