/*
 * Header file for the main_controller module.
 */

`ifndef _MAIN_CONTROLLER_H_
`define _MAIN_CONTROLLER_H_ 1

`include "main_controller/rtl/main_controller.v" // Main module include 

`endif