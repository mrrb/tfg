/*
 *
 * List of common baudrates with theirs optimal counter values [60MHz]
 *
 */

`define B921600 66
`define B460800 131
`define B256000 235
`define B230400 261
`define B153600 391
`define B128000 469

`define B115200 521
`define B57600  1042
`define B56000  1072
`define B38400  1563
`define B28800  2084
`define B19200  3125
`define B14400  4167
`define B9600   6250
`define B4800   12500
`define B2400   25000
`define B1200   50000
`define B600    100000
`define B300    200000
`define B110    545455
