/*
 * Header file for the clk_baud_pulse module.
 */

`ifndef _CLK_BAUD_PULSE_H_
`define _CLK_BAUD_PULSE_H_ 1

`include "clk_baud_pulse/rtl/clk_baud_pulse.v" // Main module include 

`endif