/*
 * Header file for the UART_Rx module.
 */

`ifndef _UART_RX_H_
`define _UART_RX_H_ 1

`include "UART/rtl/UART_Rx.v" // Main module include 

`endif