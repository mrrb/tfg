/*
 * Header file for the clk_pulse module.
 */

`ifndef _CLK_PULSE_H_
`define _CLK_PULSE_H_ 1

`include "clk_pulse/rtl/clk_pulse.v" // Main module include 

`endif