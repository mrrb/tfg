/*
 * 
 * This is the top file for the USB3300 sniffer, where all the controllers and modules are loaded
 * 
 * Modules initialization:
 *  - PLL. Module that generates the Master clock (≅100.5MHz).
 *  - UART. Module that manages the serial communication between the FPGA and the processing unit (a computer in this case).
 *  - ULPI. Module that manages the ULPI interface between the USB3300 ic and the FPGA.
 * 
 */

`default_nettype none

`define ASYNC_RESET

`ifdef ASYNC_RESET
    `define TOP_ASYNC_RESET or negedge rst
`else
    `define TOP_ASYNC_RESET
`endif

`include "./rtl/bauds.vh"

`include "./modules/UART.vh"
`include "./modules/ULPI.vh"
// `include "./modules/ULPI_WRAPPER.vh"
`include "./modules/clk_div.vh"
`include "./modules/ULPI_op_stack.vh"
`include "./modules/btn_debouncer.vh"
`include "./modules/main_controller.vh"
`include "./modules/signal_trigger.vh"

 module USB3300_sniffer #(
                          parameter DIV_TIMERS = 24,
                          parameter DIV_DEBOUNCE = 19,
                        //   parameter COUNTER_BAUDRATE = `B115200
                        //   parameter COUNTER_BAUDRATE = `B921600
                          parameter COUNTER_BAUDRATE = 16 /* Max tested baudrate 3750000 bauds -> 16 */
                         )
                         (
                          // System signals
                          input  wire clk_ice,        // 12MHz clock located in the ICEstick board
                          input  wire clk_ULPI,       // 60MHz clock from the usb3300 module

                          // ULPI signals
                          input  wire ULPI_DIR,       // ULPI DIRECTION
                          input  wire ULPI_NXT,       // ULPI NEXT
                          inout  wire [7:0]ULPI_DATA, // ULPI 8-bit parallel data
                          output wire ULPI_STP,       // ULPI STOP
                          output wire ULPI_RST,       // USB3300 RESET pin

                          // UART signals
                          input  wire UART_Rx,        // Serial Read
                          output wire UART_Tx,        // Serial Write

                          // I/O
                          input  wire [1:0]IO_BTNs,   // 
                          output wire [4:0]IO_LEDs,   // 4 (red) + 1 (green) LED's on the ICEstick board
                          output wire [2:0]IO_test
                         );

/// Config
    parameter LED_CLK_ULPI_DIV_EN = 1'b1;
    parameter LED_CLK_ICE_DIV_EN  = 1'b1;
/// End of Config

/// Reset
    wire rst;
    assign rst = btn1_debounce;
/// End of reset

/// Buttons
    wire btn1_debounce, btn2_debounce;
    wire btn2_pulse;

    btn_debouncer btn1 (
                        // System signals
                        .clk(clk_debounce),     // [Input]
                        
                        // Button
                        .btn_in(IO_BTNs[0]),    // [Input]
                        .btn_out(btn1_debounce) // [Output]
                       );

    btn_debouncer btn2 (
                        // System signals
                        .clk(clk_debounce),     // [Input]
                        
                        // Button
                        .btn_in(!IO_BTNs[1]),   // [Input]
                        .btn_out(btn2_debounce) // [Output]
                       );

    signal_trigger btn2_trigger (
                                 .clk(clk_ULPI),               // [Input]
                                 .input_signal(btn2_debounce), // [Input]
                                 .output_signal(btn2_pulse)    // [Output]
                                );
/// End of Buttons

/// Timers & clocks
    wire clk_div_ice, clk_div_ice_pulse;
    clk_div       #(.DIVIDER(DIV_TIMERS))
    clk_div_ice_m  (
                    // Clock signals
                    .clk_in(clk_ice),              // [Input]
                    .clk_out(clk_div_ice),         // [Output]
                    .clk_pulse(clk_div_ice_pulse), // [Output]

                    // Control signals
                    .enable(LED_CLK_ICE_DIV_EN)    // [Input]
                   );

    wire clk_div_ULPI, clk_div_ULPI_pulse;
    clk_div        #(.DIVIDER(DIV_TIMERS))
    clk_div_ULPI_m  (
                     // Clock signals
                     .clk_in(clk_ULPI),              // [Input]
                     .clk_out(clk_div_ULPI),         // [Output]
                     .clk_pulse(clk_div_ULPI_pulse), // [Output]

                     // Control signals
                     .enable(LED_CLK_ULPI_DIV_EN)    // [Input]
                    );

    wire clk_debounce;
    clk_div     #(.DIVIDER(DIV_DEBOUNCE))
    clk_div_btn  (
                  // Clock signals
                  .clk_in(clk_ice),       // [Input]
                  .clk_out(clk_debounce), // [Output]

                  // Control signals
                  .enable(1'b1)           // [Input]
                 );
/// End of Timers & clocks


/// Assings
    /// IO_LEDs assigns
    assign IO_LEDs[0] = clk_div_ice;   // Middle LED
    assign IO_LEDs[1] = clk_div_ULPI;  // Top LED (near FPGA ic)
    assign IO_LEDs[2] = rst;           // Left LED
    assign IO_LEDs[3] = ULPI_DIR;      // Bottom LED
    assign IO_LEDs[4] = btn2_debounce; // Right LED
/// End of Assings


/// Test assigns
    assign IO_test[0] = UART_Rx;
    assign IO_test[1] = UART_Tx;
    assign IO_test[2] = UART_send;
    // assign UART_DATA_in = UTMI_data_in_o;
    // assign UART_send    = !UART_Rx_EMPTY;
    // assign UART_NxT     = !UART_Rx_EMPTY;

    // assign UART_DATA_in = ULPI_DATA_out;
    // assign UART_DATA_in = ULPI_REG_VAL_R;
    // assign UART_DATA_in = {ULPI_REG_VAL_R[3:0], 1'b0, ULPI_busy, TOP_state_r};
    // assign UART_DATA_in = ULPI_RxCMD;
    // assign UART_DATA_in = {4'b0, ULPI_DIR, ULPI_status};
    // assign UART_DATA_in = ULPI_USB_DATA;
    // assign UART_DATA_in = UTMI_data_in_o;
    // assign UART_DATA_in = {1'b0, 1'b0, UTMI_rxvalid_o, UTMI_rxactive_o, UTMI_rxerror_o, 1'b0, 1'b1, 1'b1};

    // assign UART_DATA_in = UART_DATA_out;
    // assign UART_send    = !UART_Rx_EMPTY;
    // assign UART_NxT     = !UART_Rx_EMPTY;
/// End of Test assigns


/// PLL
    /*
     * PLL configuration
     *
     * This configuration was generated automatically
     * using the icepll tool from the IceStorm project.
     * Use at your own risk.
     *
     * Given input frequency:        12.000 MHz
     * Requested output frequency:  100.000 MHz
     * Achieved output frequency:   100.500 MHz
     */

    wire clk_ctrl;   // Generated PLL clock (≅100.5MHz)
    wire pll_locked; // Locked control signal

    SB_PLL40_CORE #(
		            .FEEDBACK_PATH("SIMPLE"),
		            .DIVR(4'b0000),		      // DIVR =  0
		            .DIVF(7'b1000010),	      // DIVF = 66
		            .DIVQ(3'b011),		      // DIVQ =  3
		            .FILTER_RANGE(3'b001)	  // FILTER_RANGE = 1
	               )
           pll_gen (
		            .LOCK(pll_locked),        // [Output]
		            .RESETB(1'b1),            // [Input]
		            .BYPASS(1'b0),            // [Input]
		            .REFERENCECLK(clk_ice),   // [Input]
		            .PLLOUTCORE(clk_ctrl)     // [Output]
		           );
/// End of PLL


/// UART
    wire [7:0]UART_DATA_in;
    wire [7:0]UART_DATA_out;
    wire UART_send;
    wire UART_TiP, UART_NrD;         // 
    wire UART_NxT;
    wire UART_Tx_FULL;                // Tx buffer status signals
    wire UART_Rx_FULL, UART_Rx_EMPTY; // Rx buffer status signals
    wire UART_Rx_clk, UART_Tx_clk;    // UART Rx/Tx clocks

    UART #(.BAUDS(COUNTER_BAUDRATE))
    UART  (
           // System signals
           .rst(rst),               // [Input]
           .clk(clk_ULPI),          // [Input]

           // UART signals
           .Rx(UART_Rx),            // [Input]
           .Tx(UART_Tx),            // [Output]
           .clk_Rx(UART_Rx_clk),    // [Output]
           .clk_Tx(UART_Tx_clk),    // [Output]

           // Data signals
           .I_DATA(UART_DATA_in),   // [Input]
           .O_DATA(UART_DATA_out),  // [Output]

           // Control signals
           .send_data(UART_send),   // [Input]
           .NxT(UART_NxT),          // [Input]
           .TiP(UART_TiP),          // [Output]
           .NrD(UART_NrD),          // [Output]
           .Tx_FULL(UART_Tx_FULL),  // [Output]
           .Rx_FULL(UART_Rx_FULL),  // [Output]
           .Rx_EMPTY(UART_Rx_EMPTY) // [Output]
          );
/// End of UART

/// ULPI INOUT tristate controller
    wire [7:0] ULPI_DATA_in, ULPI_DATA_out;

    // Yosys has only limited support for tri-state logic, so the tristate ULPI DATA bus must me manually initialized.
    // genvar i = 0;
    // generate
    //     for(i=0; i<8; i=i+1) begin : IO_TRI_DATA_GEN
    //         SB_IO      #(
    //                     .PIN_TYPE(6'b1010_01), // Input and Output Pin Function Tables. ICE Technology Library. Page 88.
    //                                             // [5:2] => PIN_OUTPUT_TRISTATE
    //                                             // [1:0] => PIN_INPUT
    //                     .PULLUP(1'b0)          // No pull-up
    //                     )
    //         IO_TRI_DATA (
    //                     .PACKAGE_PIN(ULPI_DATA[i]), // Physical tristate I/O wire
    //                     .OUTPUT_ENABLE(!ULPI_DIR),  // Control signal
    //                     .D_OUT_0(ULPI_DATA_out[i]), // 
    //                     .D_IN_0(ULPI_DATA_in[i])    // 
    //                     );
    //     end
    // endgenerate

    // Tristate selector (NOT COMPATIBLE WITH YOSYS!! [UPDATE 2019 -> Now is working just fine with the latest version of Yosys...])
    assign ULPI_DATA_in = ULPI_DATA;
    assign ULPI_DATA = (ULPI_DIR) ? 8'bz : ULPI_DATA_out; // When the PHY has the ownership of the bus, the FPGA must have the inputs in a HIGH impedance mode
                                                          // so there will not have any conflicts.
/// End of ULPI INOUT tristate controller

/// ULPI
    wire ULPI_PrW, ULPI_PrR;
    wire [2:0] ULPI_status;
    wire ULPI_busy;

    wire [5:0] ULPI_ADDR;
    wire [7:0] ULPI_REG_VAL_W, ULPI_REG_VAL_R;

    wire [7:0] ULPI_RxCMD;
    wire [1:0] ULPI_RxLineState, ULPI_RxVbusState;
    wire ULPI_RxActive, ULPI_RxError, ULPI_RxHostDisconnect, ULPI_RxID;

    wire ULPI_DATA_re, ULPI_INFO_re, ULPI_DATA_buff_full, ULPI_DATA_buff_empty, ULPI_INFO_buff_full, ULPI_INFO_buff_empty;
    wire  [7:0] ULPI_USB_DATA;
    wire [15:0] ULPI_USB_INFO_DATA;

    ULPI ULPI (
               // System signals
               .rst(rst),                                // [Input]
               .clk_ice(clk_ice),                        // [Input]
               .clk_ULPI(clk_ULPI),                      // [Input]
               
               // Control signals
               .PrW(ULPI_PrW),                           // [Input]
               .PrR(ULPI_PrR),                           // [Input]
               .status(ULPI_status),                     // [Output]
               .busy(ULPI_busy),                         // [Output]
               
               // Register signals
               .ADDR(ULPI_ADDR),                         // [Input]
               .REG_VAL_W(ULPI_REG_VAL_W),               // [Input]
               .REG_VAL_R(ULPI_REG_VAL_R),               // [Output]
               
               // Rx states
               .RxCMD(ULPI_RxCMD),                       // [Output]
               .RxLineState(ULPI_RxLineState),           // [Output]
               .RxVbusState(ULPI_RxVbusState),           // [Output]
               .RxActive(ULPI_RxActive),                 // [Output]
               .RxError(ULPI_RxError),                   // [Output]
               .RxHostDisconnect(ULPI_RxHostDisconnect), // [Output]
               .RxID(ULPI_RxID),                         // [Output]
               
               // Buffer control
               .DATA_re(ULPI_DATA_re),                   // [Input]
               .INFO_re(ULPI_INFO_re),                   // [Input]
               .USB_DATA(ULPI_USB_DATA),                 // [Output]
               .USB_INFO_DATA(ULPI_USB_INFO_DATA),       // [Output]
               .DATA_buff_full(ULPI_DATA_buff_full),     // [Output]
               .DATA_buff_empty(ULPI_DATA_buff_empty),   // [Output]
               .INFO_buff_full(ULPI_INFO_buff_full),     // [Output]
               .INFO_buff_empty(ULPI_INFO_buff_empty),   // [Output]
               
               // ULPI signals
               .DIR(ULPI_DIR),                           // [Input]
               .NXT(ULPI_NXT),                           // [Input]
               .DATA_in(ULPI_DATA_in),                   // [Input]
               .DATA_out(ULPI_DATA_out),                 // [Output]
               .STP(ULPI_STP),                           // [Output]
               .U_RST(ULPI_RST)                          // [Output]
              );
/// End of ULPI


/// ULPI op stack
    wire op_stack_pull;
    wire [15:0] op_stack_msg;
    wire op_stack_full, op_stack_empty;
    ULPI_op_stack ULPI_op_stack (
                                 // System signals
                                 .rst(rst),                      // [Input]
                                 .clk(clk_ULPI),                 // [Input]

                                 // UART Rx Buffer signals
                                 .UART_DATA(UART_DATA_out),      // [Input]
                                 .UART_Rx_EMPTY(UART_Rx_EMPTY),  // [Input]
                                 .UART_NxT(UART_NxT),            // [Output]

                                 // Stack control signals
                                 .op_stack_pull(op_stack_pull),  // [Input]
                                 .op_stack_msg(op_stack_msg),    // [Output]
                                 .op_stack_full(op_stack_full),  // [Output]
                                 .op_stack_empty(op_stack_empty) // [Output]
                                );
/// End of ULPI op stack


/// TOP controller
    main_controller main_controller (                        
                                     // System signals
                                     .rst(rst), // [Input]
                                     .clk(clk_ULPI), // [Input]
                                     .force_send(btn2_pulse),

                                     // Op stack
                                     .op_stack_msg(op_stack_msg), // [Input]
                                     .op_stack_empty(op_stack_empty), // [Input]
                                     .op_stack_pull(op_stack_pull), // [Output]

                                     // DATA ULPI signals
                                     .ULPI_USB_DATA(ULPI_USB_DATA), // [Input]
                                     .ULPI_USB_INFO_DATA(ULPI_USB_INFO_DATA), // [Input]
                                     .ULPI_DATA_buff_empty(ULPI_DATA_buff_empty), // [Input]
                                     .ULPI_INFO_buff_empty(ULPI_INFO_buff_empty), // [Input]
                                     .ULPI_DATA_re(ULPI_DATA_re), // [Output]
                                     .ULPI_INFO_re(ULPI_INFO_re), // [Output]

                                     // General ULPI signals
                                     .ULPI_busy(ULPI_busy), // [Input]

                                     // Register ULPI signals
                                     .ULPI_REG_VAL_R(ULPI_REG_VAL_R), // [Input]
                                     .ULPI_REG_VAL_W(ULPI_REG_VAL_W), // [Output]
                                     .ULPI_ADDR(ULPI_ADDR), // [Output]
                                     .ULPI_PrW(ULPI_PrW), // [Output]
                                     .ULPI_PrR(ULPI_PrR), // [Output]

                                     // UART
                                     .UART_Tx_FULL(UART_Tx_FULL), // [Input]
                                     .UART_Tx_DATA(UART_DATA_in), // [Output]
                                     .UART_send(UART_send) // [Output]
                                    );
/// End of TOP controller

endmodule