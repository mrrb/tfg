/*
 *
 * In this file are defined all the possible register address that can be read/write/set/clear in the main module.
 *
 */

 `define ADDR_CTRL_