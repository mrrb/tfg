/*
 * Header file for the clk_div module.
 */

`ifndef _CLK_DIV_H_
`define _CLK_DIV_H_ 1

`include "clk_div/rtl/clk_div.v" // Main module include 

`endif