/*
 * Header file for the UART module.
 */

`ifndef _UART_H_
`define _UART_H_ 1

`include "UART/rtl/UART.v" // Main module include 

`endif