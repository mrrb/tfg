/*
 * Header file for the ULPI module.
 */

`ifndef _ULPI_H_
`define _ULPI_H_ 1

`include "ULPI/rtl/ULPI.v" // Main module include 

`endif