/*
 * Header file for the SB_RAM40_4K module.
 */

`ifndef _SB_RAM40_4K_H_
`define _SB_RAM40_4K_H_ 1

`include "SB_RAM40_4K/rtl/SB_RAM40_4K.v" // Main module include 

`endif