/*
 * Header file for the shift_register module.
 */

`ifndef _SHIFT_REGISTER_H_
`define _SHIFT_REGISTER_H_ 1

`include "shift_register/rtl/shift_register.v" // Main module include 

`endif