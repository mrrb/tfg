/*
 * Header file for the delay module.
 */

`ifndef _DELAY_H_
`define _DELAY_H_ 1

`include "delay/rtl/delay.v" // Main module include 

`endif