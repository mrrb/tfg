/*
 * Header file for the clk_div_gen module.
 */

`ifndef _CLK_DIV_GEN_H_
`define _CLK_DIV_GEN_H_ 1

`include "clk_div_gen/rtl/clk_div_gen.v" // Main module include 

`endif