/*
 * Header file for the signal_trigger module.
 */

`ifndef _SIGNAL_TRIGGER_H_
`define _SIGNAL_TRIGGER_H_ 1

`include "signal_trigger/rtl/signal_trigger.v" // Main module include 

`endif