/*
 *
 * List of common baudrates with theirs optimal counter values
 *
 */

`define B921600 14
`define B460800 27
`define B256000 47
`define B230400 53
`define B153600 79
`define B128000 94

`define B115200 105
`define B57600  209
`define B56000  215
`define B38400  313
`define B28800  417
`define B19200  625
`define B14400  834
`define B9600   1250
`define B4800   2500
`define B2400   5000
`define B1200   10000
`define B600    20000
`define B300    40000
`define B110    109091
