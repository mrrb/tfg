/*
 * Header file for the FIFO_BRAM_SYNC module.
 */

`ifndef _FIFO_BRAM_SYNC_H_
`define _FIFO_BRAM_SYNC_H_ 1

`include "FIFO_BRAM_SYNC/rtl/FIFO_BRAM_SYNC.v" // Main module include 

`endif