/*
 * Header file for the ULPI_REG_READ module.
 */

`ifndef _ULPI_REG_READ_H_
`define _ULPI_REG_READ_H_ 1

`include "ULPI/rtl/ULPI_REG_READ.v" // Main module include 

`endif