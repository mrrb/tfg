/*
 * Header file for the SB_PLL40_CORE module.
 */

`ifndef _SB_PLL40_CORE_H_
`define _SB_PLL40_CORE_H_ 1

`include "SB_PLL40_CORE/rtl/SB_PLL40_CORE.v" // Main module include 

`endif