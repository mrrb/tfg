module top();

    

endmodule