/*
 * Header file for the REG_BANK module.
 */

`ifndef _REG_BANK_H_
`define _REG_BANK_H_ 1

`include "REG_BANK/rtl/REG_BANK.v" // Main module include 

`endif