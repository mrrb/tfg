/*
 * Header file for the btn_debouncer module.
 */

`ifndef _BTN_DEBOUNCER_H_
`define _BTN_DEBOUNCER_H_ 1

`include "btn_debouncer/rtl/btn_debouncer.v" // Main module include 

`endif